localparam UROM_BASE    = 32'h00000000;
localparam SRAM_BASE    = 32'h01000000;
localparam UART_BASE    = 32'h02000000;