localparam [7:0] BOOT   =   8'b00000001;
localparam [7:0] RUN    =   8'b00000010;

localparam UROM_BASE    = 32'h00000000;
localparam SRAM_BASE    = 32'h01000000;
localparam UART_BASE    = 32'h02000000;