localparam [7:0] USER     = 8'b00000001;
localparam [7:0] MACHINE  = 8'b00000010;