localparam [7:0] BOOT   =   8'b00000000;
localparam [7:0] RUN    =   8'b00000001;

localparam ROM_BASE  = 32'h00zzzzzz;
localparam RAM_BASE  = 32'h01zzzzzz;
localparam UART_BASE = 32'h02zzzzzz;
localparam RAMIO_BASE= 32'h03zzzzzz; 