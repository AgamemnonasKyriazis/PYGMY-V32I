localparam [7:0] ADD    =   8'b00000001 << 3'b000;
localparam [7:0] SUB    =   8'b00000001 << 3'b000;
localparam [7:0] XOR    =   8'b00000001 << 3'b100;
localparam [7:0] OR     =   8'b00000001 << 3'b110;
localparam [7:0] AND    =   8'b00000001 << 3'b111;
localparam [7:0] SLL    =   8'b00000001 << 3'b001;
localparam [7:0] SRL    =   8'b00000001 << 3'b101;
localparam [7:0] SRA    =   8'b00000001 << 3'b010;
localparam [7:0] SLT    =   8'b00000001 << 3'b010;
localparam [7:0] SLTU   =   8'b00000001 << 3'b011;